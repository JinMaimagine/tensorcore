//连接tensorcore与AXI的接口
module AXIadapter #(
)(
);
endmodule