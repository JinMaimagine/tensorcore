
module top #(
        parameter WIDTH = 6
) (
        input clk,
        input rst,
);

        

endmodule;
