//这个module用来将从systolic中收集的data转换并输出