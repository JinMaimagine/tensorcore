// ---------------------------------------------------------------------
// 32→16 converter  (combinational, round‑to‑nearest‑even)
// ---------------------------------------------------------------------
module fp32_to_fp16_conv (
    input  wire [31:0] fp32_i,
    output logic [15:0] fp16_o
);
    //------------------------------------------------------------------
    // 拆字段
    //------------------------------------------------------------------
    wire        sign  = fp32_i[31];
    wire [7:0]  exp32 = fp32_i[30:23];
    wire [22:0] man32 = fp32_i[22:0];

    //------------------------------------------------------------------
    // exp_adj = exp32 - 112  (8'h70 == 112)
    //------------------------------------------------------------------
    wire [7:0] exp_adj_full;
    SUB #(.W(8)) u_sub112 (
        .A   (exp32),
        .B   (8'h70),
        .S   (exp_adj_full),
        .Cout(/*unused*/)
    );
    wire [5:0] exp_adj = exp_adj_full[5:0];  // 用低 6 位即可

    //------------------------------------------------------------------
    // 舍入增量：+1 取决于  round_bit  &  (sticky|lsb)
    //------------------------------------------------------------------
    wire round_bit  = man32[12];
    wire sticky_bit = |man32[11:0];
    wire incr       = round_bit & (sticky_bit | man32[13]);

    wire [10:0] mant_pre  = {1'b0, man32[22:13]};        // 10+1 位
    wire [10:0] rnd_sum;
    wire        unused_c3;
    RCA #(.W(11)) u_add_rnd (
        .A   (mant_pre),
        .B   ({10'd0, incr}),        // 只在 LSB 位置加 1
        .Cin (1'b0),
        .S   (rnd_sum),
        .Cout(unused_c3)
    );

    //------------------------------------------------------------------
    // mantissa overflow 时 exponent +1
    //------------------------------------------------------------------
    wire [4:0] exp_bump;
    wire       unused_c4;
    RCA #(.W(5)) u_inc_exp (
        .A   (exp_adj[4:0]),
        .B   (5'b00001),
        .Cin (1'b0),
        .S   (exp_bump),
        .Cout(unused_c4)
    );

    //------------------------------------------------------------------
    // 主组合逻辑
    //------------------------------------------------------------------
    always_comb begin
        fp16_o = {sign, 15'd0};              // 缺省置 0

        // Inf / NaN pass-through --------------------------------------
        if (exp32 == 8'hFF) begin
            fp16_o = {sign, 5'h1F, 10'd0};
            if (man32 != 0) fp16_o[9] = 1'b1;   // qNaN
        end
        // 下溢（不支持 sub-norm 输出） -------------------------------
        else if (exp32 < 8'd103) begin        // 103 = 112-9
            fp16_o = {sign, 15'd0};
        end
        // 上溢 → Inf --------------------------------------------------
        else if (exp32 > 8'd142) begin        // 142 = 112+30
            fp16_o = {sign, 5'h1F, 10'd0};
        end
        // 正常数 ------------------------------------------------------
        else begin
            fp16_o = {sign, exp_adj[4:0], rnd_sum[9:0]};
            // mantissa overflow？
            if (rnd_sum[10]) begin
                fp16_o[14:10] = exp_bump;     // exp +1
                fp16_o[9:0]   = 10'd0;
            end
        end
    end
endmodule
