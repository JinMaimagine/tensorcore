`include "systolic.sv"
module tensorcore #(
    
)(
   
);
//TODO:控制寄存器,各种AXI接口,参考top.sv,转换到systolic所需要的接口
endmodule